module nand_gate(a,b,c);
input a,b;
output c;
nand (c,a,b);
endmodule
