module priority_encoder(input [3:0]d,output a,b,v);

always@(*)begin
case(v)
             
