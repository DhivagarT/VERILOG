module write_display;

initial begin

$display("HELLO");
$display("WORLD");
$write("HELLO\t");
$write("WORLD");

end
endmodule
