module decoder_casez;

    reg [2:0] in;
    reg [7:0] out;

    always @(*) begin
        casez(in)
            3'b000: out = 8'b00000001;
            3'b001: out = 8'b00000010;
            3'b010: out = 8'b00000100;
            3'b011: out = 8'b00001000;
            3'b100: out = 8'b00010000;
            3'b101: out = 8'b00100000;
            3'b110: out = 8'b01000000;
            3'b111: out = 8'b10000000;
            3'b1??: out = 8'b11110000;   
            default: out = 8'b00000000;
        endcase
    end

    initial begin
        $monitor("Time=%0t in=%b out=%b", $time, in, out);

        in = 3'b000; #5;
        in = 3'b001; #5;
        in = 3'b1z0; #5;  
        in = 3'b110; #5;
        in = 3'b1x1; #5;   
        in = 3'b111; #5;

        $finish;
    end

endmodule

