module gate_level1(input a,b,output out);

or (out,a,b);
endmodule

//assign out=a|b;
