module register()













































