module BINARY_to_EXCESS_3(x,a);
input [3:0]a;
output [3:0]x;

assign x = a + 4'b0011;
endmodule

